`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   20:50:03 01/19/2016
// Design Name:   adder
// Module Name:   C:/Users/schubertk/Documents/GitHub/MIPS-Lab/code/adder_test.v
// Project Name:  regs
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: adder
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module adder_test;

    // Inputs
    reg Ain;
    reg Bin;

    // Outputs
    wire add_out;

    // Instantiate the Unit Under Test (UUT)
    adder uut (
        .Ain(Ain), 
        .Bin(Bin), 
        .add_out(add_out)
    );

    initial begin
        // Initialize Inputs
        Ain = 0;
        Bin = 0;

        // Wait 100 ns for global reset to finish
        #100;
        
        // Add stimulus here

    end
      
endmodule

